// FIFO Data width
`define DATA_WD 8
// FIFO Address width
`define ADDR_WD 4
// FIFO Depth
`define FIFO_DP 16
  
// Write clock time period
`define SRC_CLK_PERIOD 100
// Read clock time period
`define DST_CLK_PERIOD 50

`define TB_IF_DEFAULT_SETUP_TIME 0.1
`define TB_IF_DEFAULT_HOLD_TIME 0.1

`define TB_IF_DEFAULT_RECOVERY_TIME 0.1
`define TB_IF_DEFAULT_REMOVAL_TIME 0.1